module ALU(
    input logic [31:0] a,
    input logic [31:0] b,

    input logic [2:0] ALU_control,
    output logic zero,overflow,negative,
    output logic [31:0] ALU_result

);


logic cout;
logic [31:0] sum;



endmodule

