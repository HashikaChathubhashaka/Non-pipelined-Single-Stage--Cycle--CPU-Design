module ALU(
    input logic [31:0] a,
    input logic [31:0] b,
    input logic [2:1] ALU_control,
    output logic carry,overflow,zero,negative,
    output logic [31:0] ALU_result

);

logic cout;
logic [31:0] sum;

    
    
endmodule