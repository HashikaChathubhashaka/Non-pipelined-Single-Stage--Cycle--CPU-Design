module branch_adder(
    input logic 
);



endmodule